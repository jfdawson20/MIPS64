module ExceptionHandler ( 



	); 
	
	
	
endmodule 