library verilog;
use verilog.vl_types.all;
entity mips64_tb is
end mips64_tb;
